module alu(
	input [15:0] A,B,
	input [3:0] ALU_Sel,
	output [15:0] ALU_Out,
	output CarryOut
	output Overflow
)
reg 7:0 ALU_Result;
wire [16:0] tmp
assign ALU_Out=ALU_result

